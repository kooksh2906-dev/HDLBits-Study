module top_module (
    output out
);
    wire GND;
    assign GND = 1'b0;
    assign out = GND;
    
endmodule