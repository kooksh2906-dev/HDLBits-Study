module top_module( output one );

// Insert your code here
wire VCC = 1'b1;
assign one = VCC;

endmodule
